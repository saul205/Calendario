{
    "2020": {
        "dia_semana": "miercoles",
        "convenio": 1792,
        "Enero": {
            "1": {
                "1": 0,
                "2": 8.5,
                "3": 7.0,
                "4": 0,
                "5": 0
            },
            "2": {
                "6": 0,
                "7": 8.5,
                "8": 8.5,
                "9": 8.5,
                "10": 7.0,
                "11": 0,
                "12": 0
            },
            "3": {
                "13": 8.5,
                "14": 8.5,
                "15": 8.5,
                "16": 8.5,
                "17": 7.0,
                "18": 0,
                "19": 0
            },
            "4": {
                "20": 8.5,
                "21": 8.5,
                "22": 8.5,
                "23": 8.5,
                "24": 7.0,
                "25": 0,
                "26": 0
            },
            "5": {
                "27": 8.5,
                "28": 8.5,
                "29": 0,
                "30": 8.5,
                "31": 7.0
            }
        },
        "Febrero": {
            "5": {
                "1": 0,
                "2": 0
            },
            "6": {
                "3": 8.5,
                "4": 8.5,
                "5": 8.5,
                "6": 8.5,
                "7": 7.0,
                "8": 0,
                "9": 0
            },
            "7": {
                "10": 8.5,
                "11": 8.5,
                "12": 8.5,
                "13": 8.5,
                "14": 7.0,
                "15": 0,
                "16": 0
            },
            "8": {
                "17": 8.5,
                "18": 8.5,
                "19": 8.5,
                "20": 8.5,
                "21": 7.0,
                "22": 0,
                "23": 0
            },
            "9": {
                "24": 8.5,
                "25": 8.5,
                "26": 8.5,
                "27": 8.5,
                "28": 7.0,
                "29": 0
            }
        },
        "Marzo": {
            "9": {
                "1": 0
            },
            "10": {
                "2": 8.5,
                "3": 8.5,
                "4": 8.5,
                "5": 0,
                "6": 7.0,
                "7": 0,
                "8": 0
            },
            "11": {
                "9": 8.5,
                "10": 8.5,
                "11": 8.5,
                "12": 8.5,
                "13": 7.0,
                "14": 0,
                "15": 0
            },
            "12": {
                "16": 8.5,
                "17": 8.5,
                "18": 8.5,
                "19": 8.5,
                "20": 7.0,
                "21": 0,
                "22": 0
            },
            "13": {
                "23": 8.5,
                "24": 8.5,
                "25": 8.5,
                "26": 8.5,
                "27": 7.0,
                "28": 0,
                "29": 0
            },
            "14": {
                "30": 8.5,
                "31": 8.5
            }
        },
        "Abril": {
            "14": {
                "1": 8.5,
                "2": 8.5,
                "3": 7.0,
                "4": 0,
                "5": 0
            },
            "15": {
                "6": 8.5,
                "7": 8.5,
                "8": 8.5,
                "9": 0,
                "10": 0,
                "11": 0,
                "12": 0
            },
            "16": {
                "13": 8.5,
                "14": 8.5,
                "15": 8.5,
                "16": 8.5,
                "17": 7.0,
                "18": 0,
                "19": 0
            },
            "17": {
                "20": 8.5,
                "21": 8.5,
                "22": 8.5,
                "23": 0,
                "24": 7.0,
                "25": 0,
                "26": 0
            },
            "18": {
                "27": 8.5,
                "28": 8.5,
                "29": 8.5,
                "30": 8.5
            }
        },
        "Mayo": {
            "18": {
                "1": 0,
                "2": 0,
                "3": 0
            },
            "19": {
                "4": 8.5,
                "5": 8.5,
                "6": 8.5,
                "7": 8.5,
                "8": 7.0,
                "9": 0,
                "10": 0
            },
            "20": {
                "11": 8.5,
                "12": 8.5,
                "13": 8.5,
                "14": 8.5,
                "15": 7.0,
                "16": 0,
                "17": 0
            },
            "21": {
                "18": 8.5,
                "19": 8.5,
                "20": 8.5,
                "21": 8.5,
                "22": 7.0,
                "23": 0,
                "24": 0
            },
            "22": {
                "25": 8.5,
                "26": 8.5,
                "27": 8.5,
                "28": 8.5,
                "29": 7.0,
                "30": 0,
                "31": 0
            }
        },
        "Junio": {
            "23": {
                "1": 8.5,
                "2": 8.5,
                "3": 8.5,
                "4": 8.5,
                "5": 7.0,
                "6": 0,
                "7": 0
            },
            "24": {
                "8": 8.5,
                "9": 8.5,
                "10": 8.5,
                "11": 8.5,
                "12": 7.0,
                "13": 0,
                "14": 0
            },
            "25": {
                "15": 8.5,
                "16": 8.5,
                "17": 8.5,
                "18": 8.5,
                "19": 7.0,
                "20": 0,
                "21": 0
            },
            "26": {
                "22": 8.5,
                "23": 8.5,
                "24": 8.5,
                "25": 8.5,
                "26": 7.0,
                "27": 0,
                "28": 0
            },
            "27": {
                "29": 8.5,
                "30": 8.5
            }
        },
        "Julio": {
            "27": {
                "1": 7.0,
                "2": 7.0,
                "3": 7.0,
                "4": 0,
                "5": 0
            },
            "28": {
                "6": 7.0,
                "7": 7.0,
                "8": 7.0,
                "9": 7.0,
                "10": 7.0,
                "11": 0,
                "12": 0
            },
            "29": {
                "13": 7.0,
                "14": 7.0,
                "15": 7.0,
                "16": 7.0,
                "17": 7.0,
                "18": 0,
                "19": 0
            },
            "30": {
                "20": 7.0,
                "21": 7.0,
                "22": 7.0,
                "23": 7.0,
                "24": 7.0,
                "25": 0,
                "26": 0
            },
            "31": {
                "27": 7.0,
                "28": 7.0,
                "29": 7.0,
                "30": 7.0,
                "31": 7.0
            }
        },
        "Agosto": {
            "31": {
                "1": 0,
                "2": 0
            },
            "32": {
                "3": 7.0,
                "4": 7.0,
                "5": 7.0,
                "6": 7.0,
                "7": 7.0,
                "8": 0,
                "9": 0
            },
            "33": {
                "10": 7.0,
                "11": 7.0,
                "12": 7.0,
                "13": 7.0,
                "14": 7.0,
                "15": 0,
                "16": 0
            },
            "34": {
                "17": 7.0,
                "18": 7.0,
                "19": 7.0,
                "20": 7.0,
                "21": 7.0,
                "22": 0,
                "23": 0
            },
            "35": {
                "24": 7.0,
                "25": 7.0,
                "26": 7.0,
                "27": 7.0,
                "28": 7.0,
                "29": 0,
                "30": 0
            },
            "36": {
                "31": 7.0
            }
        },
        "Septiembre": {
            "36": {
                "1": 8.5,
                "2": 8.5,
                "3": 8.5,
                "4": 7.0,
                "5": 0,
                "6": 0
            },
            "37": {
                "7": 8.5,
                "8": 8.5,
                "9": 8.5,
                "10": 8.5,
                "11": 7.0,
                "12": 0,
                "13": 0
            },
            "38": {
                "14": 8.5,
                "15": 8.5,
                "16": 8.5,
                "17": 8.5,
                "18": 7.0,
                "19": 0,
                "20": 0
            },
            "39": {
                "21": 8.5,
                "22": 8.5,
                "23": 8.5,
                "24": 8.5,
                "25": 7.0,
                "26": 0,
                "27": 0
            },
            "40": {
                "28": 8.5,
                "29": 8.5,
                "30": 8.5
            }
        },
        "Octubre": {
            "40": {
                "1": 8.5,
                "2": 7.0,
                "3": 0,
                "4": 0
            },
            "41": {
                "5": 8.5,
                "6": 8.5,
                "7": 8.5,
                "8": 8.5,
                "9": 7.0,
                "10": 0,
                "11": 0
            },
            "42": {
                "12": 0,
                "13": 8.5,
                "14": 8.5,
                "15": 8.5,
                "16": 7.0,
                "17": 0,
                "18": 0
            },
            "43": {
                "19": 8.5,
                "20": 8.5,
                "21": 8.5,
                "22": 8.5,
                "23": 7.0,
                "24": 0,
                "25": 0
            },
            "44": {
                "26": 8.5,
                "27": 8.5,
                "28": 8.5,
                "29": 8.5,
                "30": 7.0,
                "31": 0
            }
        },
        "Noviembre": {
            "44": {
                "1": 0
            },
            "45": {
                "2": 0,
                "3": 8.5,
                "4": 8.5,
                "5": 8.5,
                "6": 7.0,
                "7": 0,
                "8": 0
            },
            "46": {
                "9": 8.5,
                "10": 8.5,
                "11": 8.5,
                "12": 8.5,
                "13": 7.0,
                "14": 0,
                "15": 0
            },
            "47": {
                "16": 8.5,
                "17": 8.5,
                "18": 8.5,
                "19": 8.5,
                "20": 7.0,
                "21": 0,
                "22": 0
            },
            "48": {
                "23": 8.5,
                "24": 8.5,
                "25": 8.5,
                "26": 8.5,
                "27": 7.0,
                "28": 0,
                "29": 0
            },
            "49": {
                "30": 8.5
            }
        },
        "Diciembre": {
            "49": {
                "1": 8.5,
                "2": 8.5,
                "3": 8.5,
                "4": 7.0,
                "5": 0,
                "6": 0
            },
            "50": {
                "7": 0,
                "8": 0,
                "9": 8.5,
                "10": 8.5,
                "11": 7.0,
                "12": 0,
                "13": 0
            },
            "51": {
                "14": 8.5,
                "15": 8.5,
                "16": 8.5,
                "17": 8.5,
                "18": 7.0,
                "19": 0,
                "20": 0
            },
            "52": {
                "21": 8.5,
                "22": 8.5,
                "23": 8.5,
                "24": 0,
                "25": 0,
                "26": 0,
                "27": 0
            },
            "53": {
                "28": 8.5,
                "29": 0,
                "30": 8.5,
                "31": 0
            }
        }
    }
}